/***********************************************
#
#    Filename: timescale.sv
#
#    Author: ThirteenQ LJQ0 ljq1019395070@163.com
#    Description: ---
#    Create       : 2024-03-04 10:16:49
#    Last Modified: 2024-03-04 10:16:49
#
***********************************************/
`timescale 1ns/1ns
