/***********************************************
#
#    Filename: timescale.sv
#
#    Author: ThirteenQ LJQ0 ljq1019395070@163.com
#    Description: ---
#    Create       : 2024-03-14 18:42:55
#    Last Modified: 2024-03-14 18:42:55
#
***********************************************/
`timescale 1ns/1ns
