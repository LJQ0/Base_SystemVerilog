/***********************************************
#
#    Filename: PLL.sv
#
#    Author: ThirteenQ LJQ0 ljq1019395070@163.com
#    Description: 多路倍频分频
#    Create       : 2024-03-04 10:24:50
#    Last Modified: 2024-03-04 10:24:50
#
***********************************************/

