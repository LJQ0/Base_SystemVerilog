/***********************************************
#
#    Filename: timescale.sv
#
#    Author: ThirteenQ LJQ0 ljq1019395070@163.com
#    Description: ---
#    Create       : 2024-03-05 16:17:01
#    Last Modified: 2024-03-05 16:17:01
#
***********************************************/
`timescale 1ns/1ns
