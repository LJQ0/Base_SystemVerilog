/***********************************************
#
#    Filename: timescale.sv
#
#    Author: ThirteenQ LJQ0 ljq1019395070@163.com
#    Description: ---
#    Create       : 2024-03-04 15:07:15
#    Last Modified: 2024-03-04 15:07:15
#
***********************************************/
`timescale 1ns/1ns
