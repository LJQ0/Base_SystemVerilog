/***********************************************
#
#    Filename: timescale.sv
#
#    Author: ThirteenQ LJQ0 ljq1019395070@163.com
#    Description: ---
#    Create       : 2024-03-15 10:49:05
#    Last Modified: 2024-03-15 10:49:05
#
***********************************************/
`timescale 1ns/1ns
